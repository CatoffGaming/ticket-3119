module hello;
  initial begin
    $display("hello 3119");
    $finish;
  end
endmodule
